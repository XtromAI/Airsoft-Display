* Netlist for LM7805 Regulator, Voltage Divider, and Op-Amp Buffer

* 1. Power Source (V) - LiPo Battery
V_LIPO 1 0 DC 7.4  ; LiPo positive on Node 1, negative to Ground (0).

* 2. Voltage Regulator (X) - LM7805
* Format: XName Node_IN Node_GND Node_OUT ModelName
X_REG 1 2 3 LM7805 ; LM7805 regulator between IN (1), GND (2), and OUT (3).

* 3. Voltage Divider Resistors (R)
* R_TOP and R_BOT are unchanged, they still connect to Node 4.
R_TOP 1 4 2.7K     ; R_TOP (2.7K) connected between Node 1 and Node 4 (Divider Tap)
R_BOT 4 2 1K       ; R_BOT (1K) connected between Node 4 and Node 2 (LM7805 GND pin).

* 4. Op-Amp Buffer (X_BUF)
* A generic rail-to-rail Op-Amp (MODEL_OPAMP) is used, powered by the regulated 5V (Node 3) and Ground (Node 2/0).
* Configuration: Non-Inverting Input (+) connected to the Divider Tap (Node 4).
* Output (Node 5) connected back to the Inverting Input (-) for unity gain (buffer).
* The PICO_ADC now connects to the **buffer output** (Node 5).
* Format: XName +in -in +Vcc -Vcc Out ModelName
X_BUF 4 5 3 2 5 OPAMP_MODEL ; +in (4), -in (5), +Vcc (3), -Vcc (2), Out (5)

* 5. Ground Connections (Shorts)
R_GND_TIE 2 0 1u   ; Tie LM7805's GND pin (2) and Op-Amp's -Vcc pin to main PICO_GND (0).

* 6. Analysis Command (for simulation)
.OP                  ; Perform a DC Operating Point analysis.
.END                 ; End of the netlist file
